library ieee;
use ieee.std_logic_1164.all;

entity alu_tb is

end alu_tb;

architecture testbench of alu_tb is
begin
end architecture testbench;
