library ieee;
use ieee.std_logic_1164.all;

entity reg_tb is

end reg_tb;

architecture testbench of reg_tb is
begin
end architecture testbench;
