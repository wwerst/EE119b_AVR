library ieee;
use ieee.std_logic_1164.all;

entity mau_tb is

end mau_tb;

architecture testbench of mau_tb is
begin
end architecture testbench;
