library ieee;
use ieee.std_logic_1164.all;

entity avr_reg_tb is

end avr_reg_tb;

architecture testbench of avr_reg_tb is
begin
end architecture testbench;
